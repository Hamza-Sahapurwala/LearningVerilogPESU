module dff (input wire D, input wire clk, input wire rst, output reg Q);
  always @(posedge clk) 
    begin  
    if (rst)      Q <= 1'b0;     // Asynchronous reset to 0   
    else      Q <= D;        // Sample D on rising edge of clock
    end
endmodule
